.subckt sky130_fd_pr__reram_reram_cell TE BE
+ area_ox=0.1024e-12
+ Tfilament_0=3.3e-9
Xreram TE BE state_out temperature_out reram_cell_model area_ox='area_ox' Tfilament_0=Tfilament_0
.ends
